module moore (
    input wire clk, rst,
    input wire fim_pc, fim_ra, fim_rb, fim_rc, fim_rd, fim_ri, fim_ro, fim_re,
    output reg hab_pc, hab_rd, hab_ro, hab_rc, hab_re, hab_ri,
    output wire [1:0] state
);

// Declare state register
reg [1:0] sta;
assign state = sta;

// Declare states
parameter fetch = 0, decode = 1, execute = 2, conta = 3;

// Output depends only on the state
always @ (posedge clk or posedge rst) 
	begin
	  if (rst)
			sta <= fetch;
	  else
			case (sta)
				 fetch:
					  if (!fim_ri)
							sta <= fetch;
					  else
							sta <= decode;
				 decode:
					  if ((!fim_rd) || ((fim_rd) && (!fim_ro)))
							sta <= decode;
					  else if ((fim_rd) && (fim_ro))
							sta <= execute;
				 execute:
					  if (((!fim_rb) && (!fim_ra)) && (!fim_rc))
							sta <= execute;
					  else if ((!fim_rb && !fim_ra && fim_rc) || (!fim_rb && fim_ra) || (fim_rb))
							sta <= conta;
				 conta:
					  if (!fim_pc)
							sta <= conta;
					  else
							sta <= fetch;
			endcase
	end

	
always @ (sta) 
	begin
		case (sta)
			fetch:
				begin
					hab_ri <= 1'b1;
					hab_pc <= 1'b0;
					hab_rd <= 1'b0;
					hab_ro <= 1'b0;
					hab_rc <= 1'b0;
					hab_re <= 1'b0;
				end
			decode:
				begin
					hab_ro <= 1'b1;
					hab_rd <= 1'b1;
					hab_pc <= 1'b0;
					hab_rc <= 1'b0;
					hab_re <= 1'b0;
					hab_ri <= 1'b0;
				end
			execute:
				begin
					hab_re <= 1'b1;
					hab_pc <= 1'b0;
					hab_rd <= 1'b0;
					hab_ro <= 1'b0;
					hab_rc <= 1'b1;
					hab_ri <= 1'b0;
				end
			conta:
				begin
					hab_rc <= 1'b0;
					hab_pc <= 1'b1;
					hab_rd <= 1'b0;
					hab_ro <= 1'b0;
					hab_re <= 1'b0;
					hab_ri <= 1'b0;
				end
			default:
				begin
					hab_pc = 1'b0;
					hab_rd = 1'b0;
					hab_ro = 1'b0;
					hab_rc = 1'b0;
					hab_re = 1'b0;
					hab_ri = 1'b0;
				end	

		endcase
	end
	

endmodule
